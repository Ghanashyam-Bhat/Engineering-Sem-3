module and1(input wire a,b, output wire x, y);
assign y=a&b;
assign x=a|b;
endmodule
